    Mac OS X            	   2   �      �                                      ATTR       �   �   1                  �     com.apple.lastuseddate#PS       �   !  com.google.drivefs.item-id#S s��e    *�*#    1nvWv4NUyAggE15HNdD8e2xCdmJWxCZqa